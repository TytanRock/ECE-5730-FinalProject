
module MATRIX_CALCULATOR (
	clk_clk);	

	input		clk_clk;
endmodule
